
// This is one stage of an 8 stage pipelined multiplier that multiplies
// two 64-bit integers and returns the low 64 bits of the result.
// This is not an ideal multiplier but is sufficient to allow a faster clock
// period than straight multiplication.

`include "verilog/sys_defs.svh"

module mult_stage (
    input clock,
    reset,
    start,
    input [63:0] prev_sum,
    mplier,
    mcand,

    output logic [63:0] product_sum,
    next_mplier,
    next_mcand,
    output logic done
);

  parameter SHIFT = 64 / `MULT_STAGES;

  logic [63:0] partial_product, shifted_mplier, shifted_mcand;

  assign partial_product = mplier[SHIFT-1:0] * mcand;

  assign shifted_mplier  = {SHIFT'('b0), mplier[63:SHIFT]};
  assign shifted_mcand   = {mcand[63-SHIFT:0], SHIFT'('b0)};

  always_ff @(posedge clock) begin
    product_sum <= prev_sum + partial_product;
    next_mplier <= shifted_mplier;
    next_mcand  <= shifted_mcand;
  end

  always_ff @(posedge clock) begin
    if (reset) begin
      done <= 1'b0;
    end else begin
      done <= start;
    end
  end

endmodule
