// Simple bimodal branch predictor
