    Mac OS X            	   2   �      �                                      ATTR       �   �   <                  �   <  com.apple.quarantine q/0083;65f8835f;Safari;9C3630D1-0A9D-40F0-88FD-0C1F887BF25B 